`define BUFF_SIZE 16
`define DATA_BYTES_SIZE 4'h8
`define HEADER_VALUE 24'hF1
`define CH_NUM 1'h1