`define BUFF_SIZE 4
`define DATA_BYTES_SIZE 3'b100
`define HEADER_VALUE 24'hF1
`define CH_NUM 1'h1