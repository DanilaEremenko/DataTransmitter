`define BUFF_SIZE 8
`define DATA_BYTES_SIZE 4'b100