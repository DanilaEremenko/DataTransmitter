`define BUFF_SIZE 8
`define DATA_BYTES_SIZE 4'b1010
`define HEADER_VALUE 24'hF2
`define CH_NUM 2'h3